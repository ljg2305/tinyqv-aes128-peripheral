module aes128_rijndael_sbox (
    input  mode_t       mode_i,
    input  logic [7:0]  data_i, 
    output logic [7:0]  data_o
    );

    always_comb begin 
        case ({mode_i, data_i}) 
            {ENCRYPT,8'h00} :  data_o = 8'h63;
            {ENCRYPT,8'h01} :  data_o = 8'h7c;
            {ENCRYPT,8'h02} :  data_o = 8'h77;
            {ENCRYPT,8'h03} :  data_o = 8'h7b;
            {ENCRYPT,8'h04} :  data_o = 8'hf2;
            {ENCRYPT,8'h05} :  data_o = 8'h6b;
            {ENCRYPT,8'h06} :  data_o = 8'h6f;
            {ENCRYPT,8'h07} :  data_o = 8'hc5;
            {ENCRYPT,8'h08} :  data_o = 8'h30;
            {ENCRYPT,8'h09} :  data_o = 8'h01;
            {ENCRYPT,8'h0a} :  data_o = 8'h67;
            {ENCRYPT,8'h0b} :  data_o = 8'h2b;
            {ENCRYPT,8'h0c} :  data_o = 8'hfe;
            {ENCRYPT,8'h0d} :  data_o = 8'hd7;
            {ENCRYPT,8'h0e} :  data_o = 8'hab;
            {ENCRYPT,8'h0f} :  data_o = 8'h76;
            {ENCRYPT,8'h10} :  data_o = 8'hca;
            {ENCRYPT,8'h11} :  data_o = 8'h82;
            {ENCRYPT,8'h12} :  data_o = 8'hc9;
            {ENCRYPT,8'h13} :  data_o = 8'h7d;
            {ENCRYPT,8'h14} :  data_o = 8'hfa;
            {ENCRYPT,8'h15} :  data_o = 8'h59;
            {ENCRYPT,8'h16} :  data_o = 8'h47;
            {ENCRYPT,8'h17} :  data_o = 8'hf0;
            {ENCRYPT,8'h18} :  data_o = 8'had;
            {ENCRYPT,8'h19} :  data_o = 8'hd4;
            {ENCRYPT,8'h1a} :  data_o = 8'ha2;
            {ENCRYPT,8'h1b} :  data_o = 8'haf;
            {ENCRYPT,8'h1c} :  data_o = 8'h9c;
            {ENCRYPT,8'h1d} :  data_o = 8'ha4;
            {ENCRYPT,8'h1e} :  data_o = 8'h72;
            {ENCRYPT,8'h1f} :  data_o = 8'hc0;
            {ENCRYPT,8'h20} :  data_o = 8'hb7;
            {ENCRYPT,8'h21} :  data_o = 8'hfd;
            {ENCRYPT,8'h22} :  data_o = 8'h93;
            {ENCRYPT,8'h23} :  data_o = 8'h26;
            {ENCRYPT,8'h24} :  data_o = 8'h36;
            {ENCRYPT,8'h25} :  data_o = 8'h3f;
            {ENCRYPT,8'h26} :  data_o = 8'hf7;
            {ENCRYPT,8'h27} :  data_o = 8'hcc;
            {ENCRYPT,8'h28} :  data_o = 8'h34;
            {ENCRYPT,8'h29} :  data_o = 8'ha5;
            {ENCRYPT,8'h2a} :  data_o = 8'he5;
            {ENCRYPT,8'h2b} :  data_o = 8'hf1;
            {ENCRYPT,8'h2c} :  data_o = 8'h71;
            {ENCRYPT,8'h2d} :  data_o = 8'hd8;
            {ENCRYPT,8'h2e} :  data_o = 8'h31;
            {ENCRYPT,8'h2f} :  data_o = 8'h15;
            {ENCRYPT,8'h30} :  data_o = 8'h04;
            {ENCRYPT,8'h31} :  data_o = 8'hc7;
            {ENCRYPT,8'h32} :  data_o = 8'h23;
            {ENCRYPT,8'h33} :  data_o = 8'hc3;
            {ENCRYPT,8'h34} :  data_o = 8'h18;
            {ENCRYPT,8'h35} :  data_o = 8'h96;
            {ENCRYPT,8'h36} :  data_o = 8'h05;
            {ENCRYPT,8'h37} :  data_o = 8'h9a;
            {ENCRYPT,8'h38} :  data_o = 8'h07;
            {ENCRYPT,8'h39} :  data_o = 8'h12;
            {ENCRYPT,8'h3a} :  data_o = 8'h80;
            {ENCRYPT,8'h3b} :  data_o = 8'he2;
            {ENCRYPT,8'h3c} :  data_o = 8'heb;
            {ENCRYPT,8'h3d} :  data_o = 8'h27;
            {ENCRYPT,8'h3e} :  data_o = 8'hb2;
            {ENCRYPT,8'h3f} :  data_o = 8'h75;
            {ENCRYPT,8'h40} :  data_o = 8'h09;
            {ENCRYPT,8'h41} :  data_o = 8'h83;
            {ENCRYPT,8'h42} :  data_o = 8'h2c;
            {ENCRYPT,8'h43} :  data_o = 8'h1a;
            {ENCRYPT,8'h44} :  data_o = 8'h1b;
            {ENCRYPT,8'h45} :  data_o = 8'h6e;
            {ENCRYPT,8'h46} :  data_o = 8'h5a;
            {ENCRYPT,8'h47} :  data_o = 8'ha0;
            {ENCRYPT,8'h48} :  data_o = 8'h52;
            {ENCRYPT,8'h49} :  data_o = 8'h3b;
            {ENCRYPT,8'h4a} :  data_o = 8'hd6;
            {ENCRYPT,8'h4b} :  data_o = 8'hb3;
            {ENCRYPT,8'h4c} :  data_o = 8'h29;
            {ENCRYPT,8'h4d} :  data_o = 8'he3;
            {ENCRYPT,8'h4e} :  data_o = 8'h2f;
            {ENCRYPT,8'h4f} :  data_o = 8'h84;
            {ENCRYPT,8'h50} :  data_o = 8'h53;
            {ENCRYPT,8'h51} :  data_o = 8'hd1;
            {ENCRYPT,8'h52} :  data_o = 8'h00;
            {ENCRYPT,8'h53} :  data_o = 8'hed;
            {ENCRYPT,8'h54} :  data_o = 8'h20;
            {ENCRYPT,8'h55} :  data_o = 8'hfc;
            {ENCRYPT,8'h56} :  data_o = 8'hb1;
            {ENCRYPT,8'h57} :  data_o = 8'h5b;
            {ENCRYPT,8'h58} :  data_o = 8'h6a;
            {ENCRYPT,8'h59} :  data_o = 8'hcb;
            {ENCRYPT,8'h5a} :  data_o = 8'hbe;
            {ENCRYPT,8'h5b} :  data_o = 8'h39;
            {ENCRYPT,8'h5c} :  data_o = 8'h4a;
            {ENCRYPT,8'h5d} :  data_o = 8'h4c;
            {ENCRYPT,8'h5e} :  data_o = 8'h58;
            {ENCRYPT,8'h5f} :  data_o = 8'hcf;
            {ENCRYPT,8'h60} :  data_o = 8'hd0;
            {ENCRYPT,8'h61} :  data_o = 8'hef;
            {ENCRYPT,8'h62} :  data_o = 8'haa;
            {ENCRYPT,8'h63} :  data_o = 8'hfb;
            {ENCRYPT,8'h64} :  data_o = 8'h43;
            {ENCRYPT,8'h65} :  data_o = 8'h4d;
            {ENCRYPT,8'h66} :  data_o = 8'h33;
            {ENCRYPT,8'h67} :  data_o = 8'h85;
            {ENCRYPT,8'h68} :  data_o = 8'h45;
            {ENCRYPT,8'h69} :  data_o = 8'hf9;
            {ENCRYPT,8'h6a} :  data_o = 8'h02;
            {ENCRYPT,8'h6b} :  data_o = 8'h7f;
            {ENCRYPT,8'h6c} :  data_o = 8'h50;
            {ENCRYPT,8'h6d} :  data_o = 8'h3c;
            {ENCRYPT,8'h6e} :  data_o = 8'h9f;
            {ENCRYPT,8'h6f} :  data_o = 8'ha8;
            {ENCRYPT,8'h70} :  data_o = 8'h51;
            {ENCRYPT,8'h71} :  data_o = 8'ha3;
            {ENCRYPT,8'h72} :  data_o = 8'h40;
            {ENCRYPT,8'h73} :  data_o = 8'h8f;
            {ENCRYPT,8'h74} :  data_o = 8'h92;
            {ENCRYPT,8'h75} :  data_o = 8'h9d;
            {ENCRYPT,8'h76} :  data_o = 8'h38;
            {ENCRYPT,8'h77} :  data_o = 8'hf5;
            {ENCRYPT,8'h78} :  data_o = 8'hbc;
            {ENCRYPT,8'h79} :  data_o = 8'hb6;
            {ENCRYPT,8'h7a} :  data_o = 8'hda;
            {ENCRYPT,8'h7b} :  data_o = 8'h21;
            {ENCRYPT,8'h7c} :  data_o = 8'h10;
            {ENCRYPT,8'h7d} :  data_o = 8'hff;
            {ENCRYPT,8'h7e} :  data_o = 8'hf3;
            {ENCRYPT,8'h7f} :  data_o = 8'hd2;
            {ENCRYPT,8'h80} :  data_o = 8'hcd;
            {ENCRYPT,8'h81} :  data_o = 8'h0c;
            {ENCRYPT,8'h82} :  data_o = 8'h13;
            {ENCRYPT,8'h83} :  data_o = 8'hec;
            {ENCRYPT,8'h84} :  data_o = 8'h5f;
            {ENCRYPT,8'h85} :  data_o = 8'h97;
            {ENCRYPT,8'h86} :  data_o = 8'h44;
            {ENCRYPT,8'h87} :  data_o = 8'h17;
            {ENCRYPT,8'h88} :  data_o = 8'hc4;
            {ENCRYPT,8'h89} :  data_o = 8'ha7;
            {ENCRYPT,8'h8a} :  data_o = 8'h7e;
            {ENCRYPT,8'h8b} :  data_o = 8'h3d;
            {ENCRYPT,8'h8c} :  data_o = 8'h64;
            {ENCRYPT,8'h8d} :  data_o = 8'h5d;
            {ENCRYPT,8'h8e} :  data_o = 8'h19;
            {ENCRYPT,8'h8f} :  data_o = 8'h73;
            {ENCRYPT,8'h90} :  data_o = 8'h60;
            {ENCRYPT,8'h91} :  data_o = 8'h81;
            {ENCRYPT,8'h92} :  data_o = 8'h4f;
            {ENCRYPT,8'h93} :  data_o = 8'hdc;
            {ENCRYPT,8'h94} :  data_o = 8'h22;
            {ENCRYPT,8'h95} :  data_o = 8'h2a;
            {ENCRYPT,8'h96} :  data_o = 8'h90;
            {ENCRYPT,8'h97} :  data_o = 8'h88;
            {ENCRYPT,8'h98} :  data_o = 8'h46;
            {ENCRYPT,8'h99} :  data_o = 8'hee;
            {ENCRYPT,8'h9a} :  data_o = 8'hb8;
            {ENCRYPT,8'h9b} :  data_o = 8'h14;
            {ENCRYPT,8'h9c} :  data_o = 8'hde;
            {ENCRYPT,8'h9d} :  data_o = 8'h5e;
            {ENCRYPT,8'h9e} :  data_o = 8'h0b;
            {ENCRYPT,8'h9f} :  data_o = 8'hdb;
            {ENCRYPT,8'ha0} :  data_o = 8'he0;
            {ENCRYPT,8'ha1} :  data_o = 8'h32;
            {ENCRYPT,8'ha2} :  data_o = 8'h3a;
            {ENCRYPT,8'ha3} :  data_o = 8'h0a;
            {ENCRYPT,8'ha4} :  data_o = 8'h49;
            {ENCRYPT,8'ha5} :  data_o = 8'h06;
            {ENCRYPT,8'ha6} :  data_o = 8'h24;
            {ENCRYPT,8'ha7} :  data_o = 8'h5c;
            {ENCRYPT,8'ha8} :  data_o = 8'hc2;
            {ENCRYPT,8'ha9} :  data_o = 8'hd3;
            {ENCRYPT,8'haa} :  data_o = 8'hac;
            {ENCRYPT,8'hab} :  data_o = 8'h62;
            {ENCRYPT,8'hac} :  data_o = 8'h91;
            {ENCRYPT,8'had} :  data_o = 8'h95;
            {ENCRYPT,8'hae} :  data_o = 8'he4;
            {ENCRYPT,8'haf} :  data_o = 8'h79;
            {ENCRYPT,8'hb0} :  data_o = 8'he7;
            {ENCRYPT,8'hb1} :  data_o = 8'hc8;
            {ENCRYPT,8'hb2} :  data_o = 8'h37;
            {ENCRYPT,8'hb3} :  data_o = 8'h6d;
            {ENCRYPT,8'hb4} :  data_o = 8'h8d;
            {ENCRYPT,8'hb5} :  data_o = 8'hd5;
            {ENCRYPT,8'hb6} :  data_o = 8'h4e;
            {ENCRYPT,8'hb7} :  data_o = 8'ha9;
            {ENCRYPT,8'hb8} :  data_o = 8'h6c;
            {ENCRYPT,8'hb9} :  data_o = 8'h56;
            {ENCRYPT,8'hba} :  data_o = 8'hf4;
            {ENCRYPT,8'hbb} :  data_o = 8'hea;
            {ENCRYPT,8'hbc} :  data_o = 8'h65;
            {ENCRYPT,8'hbd} :  data_o = 8'h7a;
            {ENCRYPT,8'hbe} :  data_o = 8'hae;
            {ENCRYPT,8'hbf} :  data_o = 8'h08;
            {ENCRYPT,8'hc0} :  data_o = 8'hba;
            {ENCRYPT,8'hc1} :  data_o = 8'h78;
            {ENCRYPT,8'hc2} :  data_o = 8'h25;
            {ENCRYPT,8'hc3} :  data_o = 8'h2e;
            {ENCRYPT,8'hc4} :  data_o = 8'h1c;
            {ENCRYPT,8'hc5} :  data_o = 8'ha6;
            {ENCRYPT,8'hc6} :  data_o = 8'hb4;
            {ENCRYPT,8'hc7} :  data_o = 8'hc6;
            {ENCRYPT,8'hc8} :  data_o = 8'he8;
            {ENCRYPT,8'hc9} :  data_o = 8'hdd;
            {ENCRYPT,8'hca} :  data_o = 8'h74;
            {ENCRYPT,8'hcb} :  data_o = 8'h1f;
            {ENCRYPT,8'hcc} :  data_o = 8'h4b;
            {ENCRYPT,8'hcd} :  data_o = 8'hbd;
            {ENCRYPT,8'hce} :  data_o = 8'h8b;
            {ENCRYPT,8'hcf} :  data_o = 8'h8a;
            {ENCRYPT,8'hd0} :  data_o = 8'h70;
            {ENCRYPT,8'hd1} :  data_o = 8'h3e;
            {ENCRYPT,8'hd2} :  data_o = 8'hb5;
            {ENCRYPT,8'hd3} :  data_o = 8'h66;
            {ENCRYPT,8'hd4} :  data_o = 8'h48;
            {ENCRYPT,8'hd5} :  data_o = 8'h03;
            {ENCRYPT,8'hd6} :  data_o = 8'hf6;
            {ENCRYPT,8'hd7} :  data_o = 8'h0e;
            {ENCRYPT,8'hd8} :  data_o = 8'h61;
            {ENCRYPT,8'hd9} :  data_o = 8'h35;
            {ENCRYPT,8'hda} :  data_o = 8'h57;
            {ENCRYPT,8'hdb} :  data_o = 8'hb9;
            {ENCRYPT,8'hdc} :  data_o = 8'h86;
            {ENCRYPT,8'hdd} :  data_o = 8'hc1;
            {ENCRYPT,8'hde} :  data_o = 8'h1d;
            {ENCRYPT,8'hdf} :  data_o = 8'h9e;
            {ENCRYPT,8'he0} :  data_o = 8'he1;
            {ENCRYPT,8'he1} :  data_o = 8'hf8;
            {ENCRYPT,8'he2} :  data_o = 8'h98;
            {ENCRYPT,8'he3} :  data_o = 8'h11;
            {ENCRYPT,8'he4} :  data_o = 8'h69;
            {ENCRYPT,8'he5} :  data_o = 8'hd9;
            {ENCRYPT,8'he6} :  data_o = 8'h8e;
            {ENCRYPT,8'he7} :  data_o = 8'h94;
            {ENCRYPT,8'he8} :  data_o = 8'h9b;
            {ENCRYPT,8'he9} :  data_o = 8'h1e;
            {ENCRYPT,8'hea} :  data_o = 8'h87;
            {ENCRYPT,8'heb} :  data_o = 8'he9;
            {ENCRYPT,8'hec} :  data_o = 8'hce;
            {ENCRYPT,8'hed} :  data_o = 8'h55;
            {ENCRYPT,8'hee} :  data_o = 8'h28;
            {ENCRYPT,8'hef} :  data_o = 8'hdf;
            {ENCRYPT,8'hf0} :  data_o = 8'h8c;
            {ENCRYPT,8'hf1} :  data_o = 8'ha1;
            {ENCRYPT,8'hf2} :  data_o = 8'h89;
            {ENCRYPT,8'hf3} :  data_o = 8'h0d;
            {ENCRYPT,8'hf4} :  data_o = 8'hbf;
            {ENCRYPT,8'hf5} :  data_o = 8'he6;
            {ENCRYPT,8'hf6} :  data_o = 8'h42;
            {ENCRYPT,8'hf7} :  data_o = 8'h68;
            {ENCRYPT,8'hf8} :  data_o = 8'h41;
            {ENCRYPT,8'hf9} :  data_o = 8'h99;
            {ENCRYPT,8'hfa} :  data_o = 8'h2d;
            {ENCRYPT,8'hfb} :  data_o = 8'h0f;
            {ENCRYPT,8'hfc} :  data_o = 8'hb0;
            {ENCRYPT,8'hfd} :  data_o = 8'h54;
            {ENCRYPT,8'hfe} :  data_o = 8'hbb;
            {ENCRYPT,8'hff} :  data_o = 8'h16;
            {DECRYPT,8'h63} :  data_o = 8'h00;
            {DECRYPT,8'h7c} :  data_o = 8'h01;
            {DECRYPT,8'h77} :  data_o = 8'h02;
            {DECRYPT,8'h7b} :  data_o = 8'h03;
            {DECRYPT,8'hf2} :  data_o = 8'h04;
            {DECRYPT,8'h6b} :  data_o = 8'h05;
            {DECRYPT,8'h6f} :  data_o = 8'h06;
            {DECRYPT,8'hc5} :  data_o = 8'h07;
            {DECRYPT,8'h30} :  data_o = 8'h08;
            {DECRYPT,8'h01} :  data_o = 8'h09;
            {DECRYPT,8'h67} :  data_o = 8'h0a;
            {DECRYPT,8'h2b} :  data_o = 8'h0b;
            {DECRYPT,8'hfe} :  data_o = 8'h0c;
            {DECRYPT,8'hd7} :  data_o = 8'h0d;
            {DECRYPT,8'hab} :  data_o = 8'h0e;
            {DECRYPT,8'h76} :  data_o = 8'h0f;
            {DECRYPT,8'hca} :  data_o = 8'h10;
            {DECRYPT,8'h82} :  data_o = 8'h11;
            {DECRYPT,8'hc9} :  data_o = 8'h12;
            {DECRYPT,8'h7d} :  data_o = 8'h13;
            {DECRYPT,8'hfa} :  data_o = 8'h14;
            {DECRYPT,8'h59} :  data_o = 8'h15;
            {DECRYPT,8'h47} :  data_o = 8'h16;
            {DECRYPT,8'hf0} :  data_o = 8'h17;
            {DECRYPT,8'had} :  data_o = 8'h18;
            {DECRYPT,8'hd4} :  data_o = 8'h19;
            {DECRYPT,8'ha2} :  data_o = 8'h1a;
            {DECRYPT,8'haf} :  data_o = 8'h1b;
            {DECRYPT,8'h9c} :  data_o = 8'h1c;
            {DECRYPT,8'ha4} :  data_o = 8'h1d;
            {DECRYPT,8'h72} :  data_o = 8'h1e;
            {DECRYPT,8'hc0} :  data_o = 8'h1f;
            {DECRYPT,8'hb7} :  data_o = 8'h20;
            {DECRYPT,8'hfd} :  data_o = 8'h21;
            {DECRYPT,8'h93} :  data_o = 8'h22;
            {DECRYPT,8'h26} :  data_o = 8'h23;
            {DECRYPT,8'h36} :  data_o = 8'h24;
            {DECRYPT,8'h3f} :  data_o = 8'h25;
            {DECRYPT,8'hf7} :  data_o = 8'h26;
            {DECRYPT,8'hcc} :  data_o = 8'h27;
            {DECRYPT,8'h34} :  data_o = 8'h28;
            {DECRYPT,8'ha5} :  data_o = 8'h29;
            {DECRYPT,8'he5} :  data_o = 8'h2a;
            {DECRYPT,8'hf1} :  data_o = 8'h2b;
            {DECRYPT,8'h71} :  data_o = 8'h2c;
            {DECRYPT,8'hd8} :  data_o = 8'h2d;
            {DECRYPT,8'h31} :  data_o = 8'h2e;
            {DECRYPT,8'h15} :  data_o = 8'h2f;
            {DECRYPT,8'h04} :  data_o = 8'h30;
            {DECRYPT,8'hc7} :  data_o = 8'h31;
            {DECRYPT,8'h23} :  data_o = 8'h32;
            {DECRYPT,8'hc3} :  data_o = 8'h33;
            {DECRYPT,8'h18} :  data_o = 8'h34;
            {DECRYPT,8'h96} :  data_o = 8'h35;
            {DECRYPT,8'h05} :  data_o = 8'h36;
            {DECRYPT,8'h9a} :  data_o = 8'h37;
            {DECRYPT,8'h07} :  data_o = 8'h38;
            {DECRYPT,8'h12} :  data_o = 8'h39;
            {DECRYPT,8'h80} :  data_o = 8'h3a;
            {DECRYPT,8'he2} :  data_o = 8'h3b;
            {DECRYPT,8'heb} :  data_o = 8'h3c;
            {DECRYPT,8'h27} :  data_o = 8'h3d;
            {DECRYPT,8'hb2} :  data_o = 8'h3e;
            {DECRYPT,8'h75} :  data_o = 8'h3f;
            {DECRYPT,8'h09} :  data_o = 8'h40;
            {DECRYPT,8'h83} :  data_o = 8'h41;
            {DECRYPT,8'h2c} :  data_o = 8'h42;
            {DECRYPT,8'h1a} :  data_o = 8'h43;
            {DECRYPT,8'h1b} :  data_o = 8'h44;
            {DECRYPT,8'h6e} :  data_o = 8'h45;
            {DECRYPT,8'h5a} :  data_o = 8'h46;
            {DECRYPT,8'ha0} :  data_o = 8'h47;
            {DECRYPT,8'h52} :  data_o = 8'h48;
            {DECRYPT,8'h3b} :  data_o = 8'h49;
            {DECRYPT,8'hd6} :  data_o = 8'h4a;
            {DECRYPT,8'hb3} :  data_o = 8'h4b;
            {DECRYPT,8'h29} :  data_o = 8'h4c;
            {DECRYPT,8'he3} :  data_o = 8'h4d;
            {DECRYPT,8'h2f} :  data_o = 8'h4e;
            {DECRYPT,8'h84} :  data_o = 8'h4f;
            {DECRYPT,8'h53} :  data_o = 8'h50;
            {DECRYPT,8'hd1} :  data_o = 8'h51;
            {DECRYPT,8'h00} :  data_o = 8'h52;
            {DECRYPT,8'hed} :  data_o = 8'h53;
            {DECRYPT,8'h20} :  data_o = 8'h54;
            {DECRYPT,8'hfc} :  data_o = 8'h55;
            {DECRYPT,8'hb1} :  data_o = 8'h56;
            {DECRYPT,8'h5b} :  data_o = 8'h57;
            {DECRYPT,8'h6a} :  data_o = 8'h58;
            {DECRYPT,8'hcb} :  data_o = 8'h59;
            {DECRYPT,8'hbe} :  data_o = 8'h5a;
            {DECRYPT,8'h39} :  data_o = 8'h5b;
            {DECRYPT,8'h4a} :  data_o = 8'h5c;
            {DECRYPT,8'h4c} :  data_o = 8'h5d;
            {DECRYPT,8'h58} :  data_o = 8'h5e;
            {DECRYPT,8'hcf} :  data_o = 8'h5f;
            {DECRYPT,8'hd0} :  data_o = 8'h60;
            {DECRYPT,8'hef} :  data_o = 8'h61;
            {DECRYPT,8'haa} :  data_o = 8'h62;
            {DECRYPT,8'hfb} :  data_o = 8'h63;
            {DECRYPT,8'h43} :  data_o = 8'h64;
            {DECRYPT,8'h4d} :  data_o = 8'h65;
            {DECRYPT,8'h33} :  data_o = 8'h66;
            {DECRYPT,8'h85} :  data_o = 8'h67;
            {DECRYPT,8'h45} :  data_o = 8'h68;
            {DECRYPT,8'hf9} :  data_o = 8'h69;
            {DECRYPT,8'h02} :  data_o = 8'h6a;
            {DECRYPT,8'h7f} :  data_o = 8'h6b;
            {DECRYPT,8'h50} :  data_o = 8'h6c;
            {DECRYPT,8'h3c} :  data_o = 8'h6d;
            {DECRYPT,8'h9f} :  data_o = 8'h6e;
            {DECRYPT,8'ha8} :  data_o = 8'h6f;
            {DECRYPT,8'h51} :  data_o = 8'h70;
            {DECRYPT,8'ha3} :  data_o = 8'h71;
            {DECRYPT,8'h40} :  data_o = 8'h72;
            {DECRYPT,8'h8f} :  data_o = 8'h73;
            {DECRYPT,8'h92} :  data_o = 8'h74;
            {DECRYPT,8'h9d} :  data_o = 8'h75;
            {DECRYPT,8'h38} :  data_o = 8'h76;
            {DECRYPT,8'hf5} :  data_o = 8'h77;
            {DECRYPT,8'hbc} :  data_o = 8'h78;
            {DECRYPT,8'hb6} :  data_o = 8'h79;
            {DECRYPT,8'hda} :  data_o = 8'h7a;
            {DECRYPT,8'h21} :  data_o = 8'h7b;
            {DECRYPT,8'h10} :  data_o = 8'h7c;
            {DECRYPT,8'hff} :  data_o = 8'h7d;
            {DECRYPT,8'hf3} :  data_o = 8'h7e;
            {DECRYPT,8'hd2} :  data_o = 8'h7f;
            {DECRYPT,8'hcd} :  data_o = 8'h80;
            {DECRYPT,8'h0c} :  data_o = 8'h81;
            {DECRYPT,8'h13} :  data_o = 8'h82;
            {DECRYPT,8'hec} :  data_o = 8'h83;
            {DECRYPT,8'h5f} :  data_o = 8'h84;
            {DECRYPT,8'h97} :  data_o = 8'h85;
            {DECRYPT,8'h44} :  data_o = 8'h86;
            {DECRYPT,8'h17} :  data_o = 8'h87;
            {DECRYPT,8'hc4} :  data_o = 8'h88;
            {DECRYPT,8'ha7} :  data_o = 8'h89;
            {DECRYPT,8'h7e} :  data_o = 8'h8a;
            {DECRYPT,8'h3d} :  data_o = 8'h8b;
            {DECRYPT,8'h64} :  data_o = 8'h8c;
            {DECRYPT,8'h5d} :  data_o = 8'h8d;
            {DECRYPT,8'h19} :  data_o = 8'h8e;
            {DECRYPT,8'h73} :  data_o = 8'h8f;
            {DECRYPT,8'h60} :  data_o = 8'h90;
            {DECRYPT,8'h81} :  data_o = 8'h91;
            {DECRYPT,8'h4f} :  data_o = 8'h92;
            {DECRYPT,8'hdc} :  data_o = 8'h93;
            {DECRYPT,8'h22} :  data_o = 8'h94;
            {DECRYPT,8'h2a} :  data_o = 8'h95;
            {DECRYPT,8'h90} :  data_o = 8'h96;
            {DECRYPT,8'h88} :  data_o = 8'h97;
            {DECRYPT,8'h46} :  data_o = 8'h98;
            {DECRYPT,8'hee} :  data_o = 8'h99;
            {DECRYPT,8'hb8} :  data_o = 8'h9a;
            {DECRYPT,8'h14} :  data_o = 8'h9b;
            {DECRYPT,8'hde} :  data_o = 8'h9c;
            {DECRYPT,8'h5e} :  data_o = 8'h9d;
            {DECRYPT,8'h0b} :  data_o = 8'h9e;
            {DECRYPT,8'hdb} :  data_o = 8'h9f;
            {DECRYPT,8'he0} :  data_o = 8'ha0;
            {DECRYPT,8'h32} :  data_o = 8'ha1;
            {DECRYPT,8'h3a} :  data_o = 8'ha2;
            {DECRYPT,8'h0a} :  data_o = 8'ha3;
            {DECRYPT,8'h49} :  data_o = 8'ha4;
            {DECRYPT,8'h06} :  data_o = 8'ha5;
            {DECRYPT,8'h24} :  data_o = 8'ha6;
            {DECRYPT,8'h5c} :  data_o = 8'ha7;
            {DECRYPT,8'hc2} :  data_o = 8'ha8;
            {DECRYPT,8'hd3} :  data_o = 8'ha9;
            {DECRYPT,8'hac} :  data_o = 8'haa;
            {DECRYPT,8'h62} :  data_o = 8'hab;
            {DECRYPT,8'h91} :  data_o = 8'hac;
            {DECRYPT,8'h95} :  data_o = 8'had;
            {DECRYPT,8'he4} :  data_o = 8'hae;
            {DECRYPT,8'h79} :  data_o = 8'haf;
            {DECRYPT,8'he7} :  data_o = 8'hb0;
            {DECRYPT,8'hc8} :  data_o = 8'hb1;
            {DECRYPT,8'h37} :  data_o = 8'hb2;
            {DECRYPT,8'h6d} :  data_o = 8'hb3;
            {DECRYPT,8'h8d} :  data_o = 8'hb4;
            {DECRYPT,8'hd5} :  data_o = 8'hb5;
            {DECRYPT,8'h4e} :  data_o = 8'hb6;
            {DECRYPT,8'ha9} :  data_o = 8'hb7;
            {DECRYPT,8'h6c} :  data_o = 8'hb8;
            {DECRYPT,8'h56} :  data_o = 8'hb9;
            {DECRYPT,8'hf4} :  data_o = 8'hba;
            {DECRYPT,8'hea} :  data_o = 8'hbb;
            {DECRYPT,8'h65} :  data_o = 8'hbc;
            {DECRYPT,8'h7a} :  data_o = 8'hbd;
            {DECRYPT,8'hae} :  data_o = 8'hbe;
            {DECRYPT,8'h08} :  data_o = 8'hbf;
            {DECRYPT,8'hba} :  data_o = 8'hc0;
            {DECRYPT,8'h78} :  data_o = 8'hc1;
            {DECRYPT,8'h25} :  data_o = 8'hc2;
            {DECRYPT,8'h2e} :  data_o = 8'hc3;
            {DECRYPT,8'h1c} :  data_o = 8'hc4;
            {DECRYPT,8'ha6} :  data_o = 8'hc5;
            {DECRYPT,8'hb4} :  data_o = 8'hc6;
            {DECRYPT,8'hc6} :  data_o = 8'hc7;
            {DECRYPT,8'he8} :  data_o = 8'hc8;
            {DECRYPT,8'hdd} :  data_o = 8'hc9;
            {DECRYPT,8'h74} :  data_o = 8'hca;
            {DECRYPT,8'h1f} :  data_o = 8'hcb;
            {DECRYPT,8'h4b} :  data_o = 8'hcc;
            {DECRYPT,8'hbd} :  data_o = 8'hcd;
            {DECRYPT,8'h8b} :  data_o = 8'hce;
            {DECRYPT,8'h8a} :  data_o = 8'hcf;
            {DECRYPT,8'h70} :  data_o = 8'hd0;
            {DECRYPT,8'h3e} :  data_o = 8'hd1;
            {DECRYPT,8'hb5} :  data_o = 8'hd2;
            {DECRYPT,8'h66} :  data_o = 8'hd3;
            {DECRYPT,8'h48} :  data_o = 8'hd4;
            {DECRYPT,8'h03} :  data_o = 8'hd5;
            {DECRYPT,8'hf6} :  data_o = 8'hd6;
            {DECRYPT,8'h0e} :  data_o = 8'hd7;
            {DECRYPT,8'h61} :  data_o = 8'hd8;
            {DECRYPT,8'h35} :  data_o = 8'hd9;
            {DECRYPT,8'h57} :  data_o = 8'hda;
            {DECRYPT,8'hb9} :  data_o = 8'hdb;
            {DECRYPT,8'h86} :  data_o = 8'hdc;
            {DECRYPT,8'hc1} :  data_o = 8'hdd;
            {DECRYPT,8'h1d} :  data_o = 8'hde;
            {DECRYPT,8'h9e} :  data_o = 8'hdf;
            {DECRYPT,8'he1} :  data_o = 8'he0;
            {DECRYPT,8'hf8} :  data_o = 8'he1;
            {DECRYPT,8'h98} :  data_o = 8'he2;
            {DECRYPT,8'h11} :  data_o = 8'he3;
            {DECRYPT,8'h69} :  data_o = 8'he4;
            {DECRYPT,8'hd9} :  data_o = 8'he5;
            {DECRYPT,8'h8e} :  data_o = 8'he6;
            {DECRYPT,8'h94} :  data_o = 8'he7;
            {DECRYPT,8'h9b} :  data_o = 8'he8;
            {DECRYPT,8'h1e} :  data_o = 8'he9;
            {DECRYPT,8'h87} :  data_o = 8'hea;
            {DECRYPT,8'he9} :  data_o = 8'heb;
            {DECRYPT,8'hce} :  data_o = 8'hec;
            {DECRYPT,8'h55} :  data_o = 8'hed;
            {DECRYPT,8'h28} :  data_o = 8'hee;
            {DECRYPT,8'hdf} :  data_o = 8'hef;
            {DECRYPT,8'h8c} :  data_o = 8'hf0;
            {DECRYPT,8'ha1} :  data_o = 8'hf1;
            {DECRYPT,8'h89} :  data_o = 8'hf2;
            {DECRYPT,8'h0d} :  data_o = 8'hf3;
            {DECRYPT,8'hbf} :  data_o = 8'hf4;
            {DECRYPT,8'he6} :  data_o = 8'hf5;
            {DECRYPT,8'h42} :  data_o = 8'hf6;
            {DECRYPT,8'h68} :  data_o = 8'hf7;
            {DECRYPT,8'h41} :  data_o = 8'hf8;
            {DECRYPT,8'h99} :  data_o = 8'hf9;
            {DECRYPT,8'h2d} :  data_o = 8'hfa;
            {DECRYPT,8'h0f} :  data_o = 8'hfb;
            {DECRYPT,8'hb0} :  data_o = 8'hfc;
            {DECRYPT,8'h54} :  data_o = 8'hfd;
            {DECRYPT,8'hbb} :  data_o = 8'hfe;
            {DECRYPT,8'h16} :  data_o = 8'hff;
            default: data_o = 8'h00;
        endcase
    end 

endmodule 
