package aes128_type_pkg;

    typedef enum logic { ENCRYPT, DECRYPT } mode_t;

endpackage
